module all_gates(AND,OR,NOTA,NOTB,NAND,NOR,XOR,XNOR,A,B);
  input A,B;
  output AND,OR,NOTA,NOTB,NAND,NOR,XOR,XNOR;
  and(AND,A,B);
  or(OR,A,B);
  not (NOTA,A);
  not (NOTB,B);
  nand(NAND,A,B);
  nor(NOR,A,B);
  xor(XOR,A,B);
  xnor(XNOR,A,B);
endmodule
